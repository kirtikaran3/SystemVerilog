library verilog;
use verilog.vl_types.all;
entity classFunPass is
    port(
        \in\            : in     vl_logic_vector(3 downto 0)
    );
end classFunPass;
