module test(in,out); 
  
  input in; 
  output out; 
  
  assign out = in;
  
endmodule
