library verilog;
use verilog.vl_types.all;
entity classTb is
end classTb;
