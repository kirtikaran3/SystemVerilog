library verilog;
use verilog.vl_types.all;
entity dynArrTB is
end dynArrTB;
