library verilog;
use verilog.vl_types.all;
entity classFun_sv_unit is
end classFun_sv_unit;
