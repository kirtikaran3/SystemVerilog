library verilog;
use verilog.vl_types.all;
entity dynQueTB is
end dynQueTB;
